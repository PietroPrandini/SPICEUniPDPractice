* Differential Amplifier
********************************************************************************
* 3st Exercise - Fundamentals Of Electronics - a.a. 2018-2019 - UniPD - Italy  *
*                        Pietro Prandini - mat. 1097752                        *
*                                                                              *
* This work is licensed under the Creative Commons Attribution-ShareAlike 4.0  *
* International License. To view a copy of this license, visit                 *
* http://creativecommons.org/licenses/by-sa/4.0/ or send a letter to Creative  *
* Commons, PO Box 1866, Mountain View, CA 94042, USA.                          *
********************************************************************************

* Parameters
.param Vt = 0.5V
.param unCox = 200u
.param lambda = 0

.param W12 = 1.25u
.param L12 = 0.25u

.param W34 = 4.00u
.param L34 = 0.20u

.param RD = 20k

* NMOS model
.model NMOS NMOS VT0 = Vt KP = unCox LAMBDA = lambda

* Resistances
RD1 DDN D1  {RD}
RD2 DDN D2  {RD}
RD4 DDN G43 {(30/1000)*1097752}

* Transistors
MQ1 D1  G1  S12 S12 NMOS W=W12 L=L12
MQ2 S12 G2  D2  D2  NMOS W=W12 L=L12
MQ3 S12 G43 SSN SSN NMOS W=W34 L=L34
MQ4 SSN G43 G43 G43 NMOS W=W34 L=L34

* Voltage sources
VDD DDN 0 +3
VSS SSN 0 -3

* Initial conditions
.ic V(G1) = 0
.ic V(G2) = 0

* Analysis
.op

.END
