* Differential Amplifier - Differential signals
********************************************************************************
* 3st Exercise - Fundamentals Of Electronics - a.a. 2018-2019 - UniPD - Italy  *
*                        Pietro Prandini - mat. 1097752                        *
*                                                                              *
* This work is licensed under the Creative Commons Attribution-ShareAlike 4.0  *
* International License. To view a copy of this license, visit                 *
* http://creativecommons.org/licenses/by-sa/4.0/ or send a letter to Creative  *
* Commons, PO Box 1866, Mountain View, CA 94042, USA.                          *
********************************************************************************

* Parameters
.param RD = 20k

* Current sources
gm*vg2sa D2 SA G2 SA 774.76u

* Resistances
RD2 D2 0 {RD}
r0/2 SA 0 {333.2k/2}

* Voltage sources
Vi2 G2 0 sine(0 10m 10k 0 0 0)

* Analysis
.TRAN 0u 250u 0 1u

.END
