* Differential Amplifier - Differential signals
********************************************************************************
* 3st Exercise - Fundamentals Of Electronics - a.a. 2018-2019 - UniPD - Italy  *
*                        Pietro Prandini - mat. 1097752                        *
*                                                                              *
* This work is licensed under the Creative Commons Attribution-ShareAlike 4.0  *
* International License. To view a copy of this license, visit                 *
* http://creativecommons.org/licenses/by-sa/4.0/ or send a letter to Creative  *
* Commons, PO Box 1866, Mountain View, CA 94042, USA.                          *
********************************************************************************

* Parameters
.param RD = 20k

* Current sources
gm*vg1s1 D1 0 G1 0 774.76u
gm*vg2s2 D2 0 G2 0 774.76u
gm*vd4ss4 D4 0 D4 0 547.80
gm*vd4ss3 SA 0 D4 0 547.80

* Resistances
RD1 0 D1 {RD}
RD2 0 D2 {RD}
RD4 0 D4 33k
r0 0 SA 333.2k

* Voltage sources
Vi1 G1 0 sine(0 10m 10k 0 0 0)
Vi2 0 G2 sine(0 10m 10k 0 0 0)

* Analysis
.TRAN 0u 250u 0 1u

.END
