* NMOS amplifier
********************************************************************************
* 2st Exercise - Fundamentals Of Electronics - a.a. 2018-2019 - UniPD - Italy  *
*                        Pietro Prandini - mat. 1097752                        *
*                                                                              *
* This work is licensed under the Creative Commons Attribution-ShareAlike 4.0  *
* International License. To view a copy of this license, visit                 *
* http://creativecommons.org/licenses/by-sa/4.0/ or send a letter to Creative  *
* Commons, PO Box 1866, Mountain View, CA 94042, USA.                          *
********************************************************************************

* NMOS model
.model NMOS NMOS VT0 = 1V KP = 4m LAMBDA = 0

* Generators
*VDD NDD 0 15V

* Resistances
RG1 VDD VG 2.19550MEG
RG2 VG 0 1097752
RD VDD VD 8K
RS VS 0 7K

* Transistors
M1 VD VG VS VS NMOS

* Initial conditions
.ic V(VDD) = 15V

* Analysis
.op

.END
