* Differential Amplifier - Static conditions - Differential Amplifier part
********************************************************************************
* 3st Exercise - Fundamentals Of Electronics - a.a. 2018-2019 - UniPD - Italy  *
*                        Pietro Prandini - mat. 1097752                        *
*                                                                              *
* This work is licensed under the Creative Commons Attribution-ShareAlike 4.0  *
* International License. To view a copy of this license, visit                 *
* http://creativecommons.org/licenses/by-sa/4.0/ or send a letter to Creative  *
* Commons, PO Box 1866, Mountain View, CA 94042, USA.                          *
********************************************************************************

* Parameters
.param RD = 20k

* NMOS models
.model NA NMOS VT0=0.5 KP=200u LAMBDA=0 W=4.00u L=0.20u

* Current sources
ISA/2 SA SS {150.06433u/2}

* Resistances
RD1 DD D1 {RD}

* Transistors
M1 D1 G1 SA SA NA

* Voltage sources
VDD DD 0 3
VSS SS 0 -3
Vi1 G1 0 0

* Analysis
.op

.END
