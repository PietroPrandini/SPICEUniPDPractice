* Differential Amplifier
********************************************************************************
* 3st Exercise - Fundamentals Of Electronics - a.a. 2018-2019 - UniPD - Italy  *
*                        Pietro Prandini - mat. 1097752                        *
*                                                                              *
* This work is licensed under the Creative Commons Attribution-ShareAlike 4.0  *
* International License. To view a copy of this license, visit                 *
* http://creativecommons.org/licenses/by-sa/4.0/ or send a letter to Creative  *
* Commons, PO Box 1866, Mountain View, CA 94042, USA.                          *
********************************************************************************

* Parameters
.param RD = 20k

.param VG1 = 0
.param VG2 = 0

* NMOS model
*.model ND NMOS VT0=0.5 KP=200u LAMBDA=0 W=4.00u L=0.20u
.model NMOS NMOS VT0=0.5 KP=200u LAMBDA=0

* Resistances
*RD1 DD D1 {RD}
*RD2 DD D2 {RD}
RD4 DD D4 33k

* Transistors
*M1 D1 G1 SA SA ND
*M2 SA G2 D2 D2 ND
*M3 SA D4 SS SS NS
M4 D4 D4 SS SS NMOS  W=1.25u L=0.25u

* Voltage sources
VDD DD 0 3
VSS 0 SS 3
*Vi1 G1 0 {VG1}
*Vi2 G2 0 {VG2}

* Analysis
.op

.END
